-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Sun Nov 17 20:43:11 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY \4b_2to1MUX\ IS 
	PORT
	(
		S :  IN  STD_LOGIC;
		I0 :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		I1 :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		F :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END \4b_2to1MUX\;

ARCHITECTURE bdf_type OF \4b_2to1MUX\ IS 

COMPONENT \2to1mux\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 S : IN STD_LOGIC;
		 F : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	F_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN 



b2v_inst : \2to1mux\
PORT MAP(A => I0(0),
		 B => I1(0),
		 S => S,
		 F => F_ALTERA_SYNTHESIZED(0));


b2v_inst1 : \2to1mux\
PORT MAP(A => I0(1),
		 B => I1(1),
		 S => S,
		 F => F_ALTERA_SYNTHESIZED(1));


b2v_inst2 : \2to1mux\
PORT MAP(A => I0(2),
		 B => I1(2),
		 S => S,
		 F => F_ALTERA_SYNTHESIZED(2));


b2v_inst3 : \2to1mux\
PORT MAP(A => I0(3),
		 B => I1(3),
		 S => S,
		 F => F_ALTERA_SYNTHESIZED(3));

F <= F_ALTERA_SYNTHESIZED;

END bdf_type;